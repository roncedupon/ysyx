module EXU(
    input clk,
    input rst
);
endmodule