module top(
	    input clk,
	        input rst_n,
		    output clk_o,
		        output rst_n_o
		);
		assign clk_o=clk;
		assign rst_n_o=rst_n;
		endmodule
