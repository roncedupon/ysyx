module adder(input a,input b,output c);
endmodule