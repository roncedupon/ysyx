module IDU(

);
endmodule