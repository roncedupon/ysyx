module IFU(//取指单元
    input clk,//输入时钟

);
endmodule
